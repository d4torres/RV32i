`define RISCV_FORMAL
`define NRET 1
`define XLEN 32
`define ILEN 32
`define DEBUG