`define RISCV_FORMAL
`define DEBUG
